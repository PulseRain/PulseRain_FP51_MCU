// Altera_unique_chip_ID.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module Altera_unique_chip_ID (
		input  wire        clkin,      //  clkin.clk
		input  wire        reset,      //  reset.reset
		output wire        data_valid, // output.valid
		output wire [63:0] chip_id     //       .data
	);

	altchip_id #(
		.DEVICE_FAMILY ("MAX 10"),
		.ID_VALUE      (64'b0001001000110100010101100111100010101010101110111100110011011101),
		.ID_VALUE_STR  ("00000000aabbccdd")
	) altera_unique_chip_id_inst (
		.clkin      (clkin),      //  clkin.clk
		.reset      (reset),      //  reset.reset
		.data_valid (data_valid), // output.valid
		.chip_id    (chip_id)     //       .data
	);

endmodule
